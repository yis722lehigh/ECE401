module ROM(out,address);
	output reg [31:0] out;
	input [31:0] address; 
	//input clock;
	always @(address) begin
		case (address)
		
		   /*32'd00: out = 32'h00000000;
			32'd04: out = 32'h00400513;//addi x10,x0,4   0000 0000 0100 0101 0000 0101 0001 0011
			32'd08: out = 32'h00100713; //addi x14,x0,1  0000 0000 0001 0000 0000 0111 0001 0011 
			
			32'd12: out = 32'h00e507b3; // add x15,x10,x14 0000 000 01110 01010 000 01111 0110011 // 0000 0000 1110 0101 0000 0111 1011 0011 //0111 1010
			32'd16: out = 32'h00178813; // addi x16,x15,1 0000 0000 0001 01111 000 10000 0010011 // 0000 0000 0001 0111 1000 1000 0001 0011*/
			
			
			32'd00: out = 32'h00000000;
			/*32'd04: out = 32'b00400513;//addi x10,x0,4   0000 0000 0100 0101 0000 0101 0001 0011
			32'd08: out = 32'b00100713; //addi x14,x0,1  0000 0000 0001 0000 0000 0111 0001 0011 
			
			32'd12: out = 32'h00e507b3; // add x15,x10,x14 0000 000 01110 01010 000 01111 0110011 // 0000 0000 1110 0101 0000 0111 1011 0011 //0111 1010
			32'd16: out = 32'h00178813; // addi x16,x15,1 0000 0000 0001 01111 000 10000 0010011 // 0000 0000 0001 0111 1000 1000 0001 0011
			
			*/                 //imm        rs1 funct3 rd   opcode
	      32'd04: out = 32'b00000000010000000000010100010011;//addi x I-- 
         32'd08: out = 32'b00000000000100000000011100010011;//addi I--
         32'd12: out = 32'b00000000111001010000011110110011; //add R--
         32'd16: out = 32'b00000000111101010010001000010011;//I--
         32'd20: out = 32'b00000000010001010010100000000011;//I--
         32'd24: out = 32'b00000000111110000000001001000111;
         32'd28: out = 32'b00000000111001010100011110110011;//R--
         32'd32: out = 32'b01000000111001010000011000110011;//R--

			
			
			
		
		
			/*32'd00: out = 32'h00450013;//addi x13,x0,4   0000 0000 0100 0101 0000 0000 0001 0011
			32'd04: out = 32'h00100713; //addi x14,x0,1  0000 0000 0001 0000 0000 0111 0001 0011 
			32'd08: out = 32'h00d707b3; // add x15,x14,x13 0000 0000 1101 0111 0000 0111 1011 0011 
			*/
			
			
			/*8'd00: out = 32'h00450693;//addi a3,a0,4   
			8'd04: out = 32'h00100713; //addi a4,x0,1 
			8'd08: out = 32'h00b76463; // bltu a4,a1,10 --Outer Loop:
			8'd12: out = 32'h00008067; //addi x0,x1,0  --Exit Outer Loop:
			8'd16: out = 32'h0006a803; //a6,0(a3) --Continue Outer Loop:
			8'd20: out = 32'h00068613; //a2,a3,0
			8'd24: out = 32'h00070793; //a5,a4,0
			8'd28: out = 32'hffc62883; //a7,-4(a2) --Inner Loop:
			8'd32: out = 32'h01185a63; //a6,a7,34
			8'd36: out = 32'h01162023; //a7,0(a2)
			8'd40: out = 32'hfff78793; //a5,a5,-1
			8'd44: out = 32'hffc60613; //a2,a2,-4
			8'd48: out = 32'hfe0796e3; //a5,x10,1c
			8'd52: out = 32'h00279793; //a5,a5,0x2 --Exit inner loop
			8'd56: out = 32'h00f507b3; //a5,a0,a5
			8'd60: out = 32'h0107a023; //a6,0(a5)
			8'd64: out = 32'h00170713; //a4,a4,1
			8'd68: out = 32'h00468693; //a3,a3,4
			8'd72: out = 32'hfc1ff06f; //x0,8*/
			
			
			
			default:  out = 32'h00000000; 
		endcase
	end
endmodule
